library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity reg14bits is 
    port(   clk, reset, wr_en : in std_logic;
            data_in : in unsigned(13 downto 0);
            data_out : out unsigned(13 downto 0)
    );
end entity;

architecture a_reg14bits of reg14bits is 
    signal registro: unsigned(13 downto 0);
begin

    process(clk, reset, wr_en)
    begin
        if reset='1' then
            registro <= "00000000000000";
        elsif wr_en='1' then
            if rising_edge(clk) then
                registro <= data_in;
            end if;
        end if;
    end process;

    data_out <= registro;
end architecture;
